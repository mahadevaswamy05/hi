
class packet;

rand bit [3:0] a;
endclass
