mahadevaswamy
27-01-2022
place:manipal
