int a;
module name;
endmodule:wq
