`define M1 50

module test;
initial begin
    $display("output M1",`M1);
  end
  endmodule

