module pkg;
`define WIDTH 20; 
  function int two(int a,b);
    int c;
    c=a+b;
    $display("the valeue a=%0d b=%0d c=%0d",a,b,c);
    return (c);
  endfunction

  endmodule

