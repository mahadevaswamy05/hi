//interface code

interface add_if();
 logic [3:0]a;
 logic [3:0]b;
 logic clk;
 logic cin;
 logic [3:0]sum;
 logic cout;
 logic rst;

endinterface 
