<<<<<<< HEAD
mahadevaswamy
27-01-2022
place:manipal
=======
int a;
module name;
endmodule:wq
>>>>>>> main
