module tb;
import pkg::*;

initial begin
  pkg::two(2,3);
end
endmodule
