just go the visual mode then ctrl+v it will selecting the letter vertically then type shift + i
and then type command (//) then esc . //this is for the multiply line commands at time.

ctrl+g for knowing the file name in the opening other file
/ searching keyword and n for going to next words
? searching the words in the backword manner

marking some location and jumping to that location
ma for making the loaction
'a for jumping to that location like a marked location 
for multiply mark locations mg for first marked locations or mk for second marked locations
'g for jumping into first maked location and 'k for second marked locations 
zz for middle of the screen

. for repeating the previous command just it will do the last command repeating 
s/p/packet for you can select the particular season and we can do the replace of the word
ctrl+v for seleting the words in the from of vertical
== for indentation
ctrl+v
d$ for where cursor is pointing to end line it will delete.
e for jumping the one word to another word
w for jumping the one word to another word
yiw for copying the particular word 
ciw for cutting the particular word
% for jumping the one statrting parentheses to ending parenthenses but cursor as to pointing to starting parentheses
%d for it will delete the inside the parentheses things parentheses

// >>
//  << 
you write this things in the file which file you wanted to do indentation  go to visual mode and then type >> for right identation << for left side indentation

