[?1049h[?1h=[1;24r[?12;25h[?12l[?25h[27m[m[38;5;252m[48;5;234m[H[2J[?25l[24;1H"dynamic_" [New File][1;1H[38;5;240m[48;5;234m  1 
~                                                                               [3;1H~                                                                               [4;1H~                                                                               [5;1H~                                                                               [6;1H~                                                                               [7;1H~                                                                               [8;1H~                                                                               [9;1H~                                                                               [10;1H~                                                                               [11;1H~                                                                               [12;1H~                                                                               [13;1H~                                                                               [14;1H~                                                                               [15;1H~                                                                               [16;1H~                                                                               [17;1H~                                                                               [18;1H~                                                                               [19;1H~                                                                               [20;1H~                                                                               [21;1H~                                                                               [22;1H~                                                                               [23;1H~                                                                               [m[38;5;252m[48;5;234m[24;63H0,0-1[9CAll[1;5H[?12l[?25h[24;1H
[39;49m[?1l>[?1049l[?1049h[?1h=[?12;25h[?12l[?25h[27m[m[38;5;252m[48;5;234m[H[2J[?25l[1;1H[38;5;240m[48;5;234m  1 
~                                                                               [3;1H~                                                                               [4;1H~                                                                               [5;1H~                                                                               [6;1H~                                                                               [7;1H~                                                                               [8;1H~                                                                               [9;1H~                                                                               [10;1H~                                                                               [11;1H~                                                                               [12;1H~                                                                               [13;1H~                                                                               [14;1H~                                                                               [15;1H~                                                                               [16;1H~                                                                               [17;1H~                                                                               [18;1H~                                                                               [19;1H~                                                                               [20;1H~                                                                               [21;1H~                                                                               [22;1H~                                                                               [23;1H~                                                                               [m[38;5;252m[48;5;234m[24;63H0,0-1[9CAll[1;5H[?12l[?25h[24;1H[39;49m[?1l>[?1049lVim: Caught deadly signal TERM
Vim: Finished.
[24;1H[27m[m[38;5;252m[48;5;234m[39;49m